module seven_segment (
input [3:0]i,
output reg [6:0]o
);


// HEX out - rewire DE2
//  ---a---
// |       |
// f       b
// |       |
//  ---g---
// |       |
// e       c
// |       |
//  ---d---
always @(*)
	begin
		case (i)	    // abcdefg
			4'b0000: o = 7'b0000001;//0
			4'b0001: o = 7'b1001111;//1
			4'b0010: o = 7'b0010010;//2
			4'b0011: o = 7'b0000110;//3
		
			4'b0100: o = 7'b1001100;//4
			4'b0101: o = 7'b0100100;//5
			4'b0110: o = 7'b0100000;//6
			4'b0111: o = 7'b0001111;//7
		
			4'b1000: o = 7'b0000000;//8
			4'b1001: o = 7'b0000100;//9
			4'b1010: o = 7'b0001000;//a
			4'b1011: o = 7'b1100000;//b
		
			4'b1100: o = 7'b0110001;//c
			4'b1101: o = 7'b1000010;//d
			4'b1110: o = 7'b0110000;//e
			4'b1111: o = 7'b0111000;//f
		
			default: o = 7'b1111111;

		endcase
	end

endmodule